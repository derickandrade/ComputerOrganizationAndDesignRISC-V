library verilog;
use verilog.vl_types.all;
entity ulaRV_vlg_vec_tst is
end ulaRV_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity ulaRISCV_vlg_vec_tst is
end ulaRISCV_vlg_vec_tst;
